/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
    // Do a multiplication to create a bunch of gates
    logic [15:0] product;
    
    always @(posedge clk, negedge rst_n) begin
        if (!rst_n) begin
            product <= '0;
        end else begin
            product <= ui_in * uio_in;
        end

    end
    
    assign uo_out  = product[7:0];
    assign uio_out = product[15:8];
    assign uio_oe  = '0;

    // List all unused inputs to prevent warnings
    wire _unused = ena;

endmodule
